`timescale 1ns/1ps
module tb_cb_seg();
reg clk, reset, wreq_tb, wreq_size;
reg [7:0] tb_in;
reg[11:0] tb_size_in;

//wire filling, crc, start, stop, cb_size;
//wire[7:0] cb_data;

wire empty_itl,empty_enc;
reg  rreq_itl, rreq_enc;

wire[9:0] q_enc;
wire size_enc, start_enc;
wire[7:0] data_enc;

wire[9:0] q_itl;
wire size_itl, start_itl;
wire[7:0] data_itl;

assign data_itl = q_itl[9:2];
assign size_itl = q_itl[1];
assign start_itl = q_itl[0];

assign data_enc = q_enc[9:2];
assign size_enc = q_enc[1];
assign start_enc = q_enc[0];


cb_seg test_obj(
    .clk(clk),
    .reset(reset),
    .tb_in(tb_in),
    .wreq_data(wreq_tb),
    .tb_size_in(tb_size_in),  
    .wreq_size(wreq_size),
	 
	 .rreq_itl_fifo(rreq_itl),
	 .q_itl_fifo(q_itl), //{data, size, start}
	 .empty_itl_fifo(empty_itl),
	 
	 //Encoder FIFO Ports
	 .rreq_enc_fifo(rreq_enc),
	 .q_enc_fifo(q_enc),  //{data, size, start, crc, filling}
	 .empty_enc_fifo(empty_enc)
	 

//    .filling(filling),
//    .crc(crc),
//    .start(start),
//    //.stop(stop),
//    .cb_size(cb_size),
//    .cb_data(cb_data) 
);


//integer length = 7024 = 8*878;
integer length = 878;
integer iterations = 925, i, k;
integer record_start= 0;
reg [7:0] check_out;
reg switch = 1'b0;

wire[7023:0] input_vector = 7024'b0101011101000011111000101001010101101111110110101010111000001011001000101001000011111100110001110001000010000110111100010010101101011110000001100101110110010110111110101001101011111001101100011101111001011100010110111100100011110100100110110011100100000111110100100000000100010100110110100100110000010011101000010111000110001101100011110001010110111111111011001110001011100010111000100111001010111101011010001100010101001101100000101001101100111111011001110110000011100011101111111010000001100010000100100100111101100001000010110101000001000111010001100011100110010000101100010101010100001010100110100100110101100001011101001001111001000001011001010001000111101100000101010010011010000010011001101101100011110011111000000000000011001100110100101010100100100010000010101111010010010111111010011000110100001101101100000100101110010010110000100110100110111110000001001011100001010000010101010001110011111110101111100101111111010111001011001010101101000111000000101111111010011101110101110000000001100011110101011011111000011001001000111100011111010001011001010111100000000100001000111110110101001001100110001100011011111111110011000101110110010110101111110100101011000110100010111111011001100100001000001101110110110110001011100110101110011001010000101011100000011001101111000010010010010001111101101110011100000001110000010101000100000000101100100000011011111100111001101000000010111101111101000001010111001111101010101011000011001010110000011010100010001011000111000111001000110001110001110110010110011100100111001100111000010001100100100101010111001110110000010100000010000010010011101001000111001001111000000010110110000101000001101100111101011100101000111011110100011010100001110000001111111101011101000111110000110110110010110010110001010001111010111001011100010010010010010011110000110101100010001101101000110001010110101100000111110001000000010010001101100110110111101011111111001000001011110100111100111110110111110100101001111000111011001011000001111111001110010111110111110110101101110000010110010010110001110001110010110010101111001100111100101100001101111010010111001101010011110111110000011111110010110110100010100111110010100100001101011101110101001001110000110111010111110111111000111100011000000011001100100111000001110001000011000011111011000101010100111011111100010111111111000101010100101010111101110101111001111010110100010000011101100101101001011111100110010010100000100001111111111011011100011000010111011101010110010100101100111000100101101000100011110010110110100011100100111111110001100001000011100101010011001100010101000101111011010110100101100111001001100100100000100110001010000101000101100000001100100100001101001001010111010010001101101000101100101100100011100000011110011010011101010001110000000011011111010111001011000011101010111100010011011001010110100100010000101011010011100000111001100111101001110010111111000101011100001010110101110000100100111001000010111100110011001001000111011011111001001011111101111010100111010101010011010010101011001000110101011111111110000111011101001100101110000000010000011100010010010101100000010100100000001110101110000101001010101010000100010101110000001011101111011001010000010000010001111110110110000111100101101110001110000000011111110110000001011111010110101111101110111110011101111000010111111110000001111110011010101010000000000010010000011001110100100110010001000100110110111110111000011110100011100101101111101010101010111001100001000011001110110001101001101101001001000110000110011001001110000100001000010000101011000011010110111000101110010101001000111000101110010000010100001010101110011110111101100011101011100001111010010101000100110101101001001010010001110011000101111011001010101101101100101001111111001101110000111101000110001010001100000010101111110110010110101111010000101001000101001100000011100101010101010101110011110100101111100011110100011010010100010110001010111000100010000011110100101010111001101000000101000011011100101000000101010011000100100110111100000001010010010110111000110001001010111100101010101010010100000011010111100111110111101100010111010010110110001000110011001100111111101111100101010110011001111110100101000111000110110100010101111100011110110011010100100010101010100101000010001100111001100000111111010001001100110111101101100110110011101100100101001100101000101100110110101001000001000101001000010000000110001110110110111000001001001100110101110101100010011110010100111101001011011110110011001101110001100111010111010101111010100001011111100110100000010011000111100111110111000101000010010010010000011000110000001110011110001111011011100111010100011110100110001111100111111001100010010100000001010100101000111110110100001101111111000000000111011111100101011110010001111110100001010000010101011010100001011011110111000011111110011001111011000010011110110010010100111110000111000010000111001100000000001111010000100110001101111111010010110010101000010110100110110110011101000000010001111001000011001101001000011011001010001011100101001111101111110011000101110111111110000111011100110010000110100011111000111000000011110001111100000100111111111111001011100100001110110110000001010100011001100001111011000011111110110010000111001001100000000110001000110000011001011101011011101101100010100101000001100111100110001111110010010001100000101000100111000100000110000100011001011010001010011111101010111111111010001011010011110001111111101101110101000001011001001000011110111100111101010101010110111001101100011101110110001010110101101110000000000010101101100011100001010011000010110101110100011010110110000000100000100001101111011011000000011110101001011010110110111000011001010011110000000100100110100100000010001110100010010101100001010100101001101110101100011011100010111101100100001001011111100101100110111000010100000001010100000010100001000111111110000010000111110100001000011000110110011001000000010001001100111101001101110000100001011001010000110111010100110001011000111100111111111000111001101101001100111110010011100001000011111001010111100010110100000101010011111110100011000001111001101100101101100100111010010010110001000000110101111010000010110000110010100010010010001011000000111001100001000001101010101111011010001010111100111011011110110111110000010001000111111111000000010001100001111010111111100001100011110111010011100001100011010100110011001111000100101000111000011100110010101011000011011000000000000010100100100011111111110001000010111100000111000100010010110100000101110011010110100101011011000111111000111011011000010001101010001010010001011111111001100001000010001110001111110101111011011101101110101111000010101100111111111001000100010100000010000010000100001011110010010100111011011010011100011100100000011011010001001011001001111010111000111100001000010110010101101110001110001001100110111110001110011100100111100110000001100100110010010101110000000011010001100100101011110101010111100111101101111100100111000100101111110001000001011101000101001001100101101101010100100100100100000001001010111011001101010111100010010010000000010000011101010010101101011110001001011100111110111001110000111100;

wire[1031:0] cb1_data = 1032'b111101101000101011110011101101111011011111000001000100011111111100000001000110000111101011111110000110001111011101001110000110001101010011001100111100010010100011100001110011001010101100001101100000000000001010010010001111111111000100001011110000011100010001001011010000010111001101011010010101101100011111100011101101100001000110101000101001000101111111100110000100001000111000111111010111101101110110111010111100001010110011111111100100010001010000001000001000010000101111001001010011101101101001110001110010000001101101000100101100100111101011100011110000100001011001010110111000111000100110011011111000111001110010011110011000000110010011001001010111000000001101000110010010101111010101011110011110110111110010011100010010111111000100000101110100010100100110010110110101010010010010010000000100101011101100110101011110001001001000000001000001110101001010110101111000100101110011111011100111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire[23:0] cb1_crc = 24'b000010110010111100011011;
//From MSB to LSB
wire[1055:0] output_vector1 = {cb1_crc, cb1_data};


wire[6119:0] cb2_data = 6120'b010101110100001111100010100101010110111111011010101011100000101100100010100100001111110011000111000100001000011011110001001010110101111000000110010111011001011011111010100110101111100110110001110111100101110001011011110010001111010010011011001110010000011111010010000000010001010011011010010011000001001110100001011100011000110110001111000101011011111111101100111000101110001011100010011100101011110101101000110001010100110110000010100110110011111101100111011000001110001110111111101000000110001000010010010011110110000100001011010100000100011101000110001110011001000010110001010101010000101010011010010011010110000101110100100111100100000101100101000100011110110000010101001001101000001001100110110110001111001111100000000000001100110011010010101010010010001000001010111101001001011111101001100011010000110110110000010010111001001011000010011010011011111000000100101110000101000001010101000111001111111010111110010111111101011100101100101010110100011100000010111111101001110111010111000000000110001111010101101111100001100100100011110001111101000101100101011110000000010000100011111011010100100110011000110001101111111111001100010111011001011010111111010010101100011010001011111101100110010000100000110111011011011000101110011010111001100101000010101110000001100110111100001001001001000111110110111001110000000111000001010100010000000010110010000001101111110011100110100000001011110111110100000101011100111110101010101100001100101011000001101010001000101100011100011100100011000111000111011001011001110010011100110011100001000110010010010101011100111011000001010000001000001001001110100100011100100111100000001011011000010100000110110011110101110010100011101111010001101010000111000000111111110101110100011111000011011011001011001011000101000111101011100101110001001001001001001111000011010110001000110110100011000101011010110000011111000100000001001000110110011011011110101111111100100000101111010011110011111011011111010010100111100011101100101100000111111100111001011111011111011010110111000001011001001011000111000111001011001010111100110011110010110000110111101001011100110101001111011111000001111111001011011010001010011111001010010000110101110111010100100111000011011101011111011111100011110001100000001100110010011100000111000100001100001111101100010101010011101111110001011111111100010101010010101011110111010111100111101011010001000001110110010110100101111110011001001010000010000111111111101101110001100001011101110101011001010010110011100010010110100010001111001011011010001110010011111111000110000100001110010101001100110001010100010111101101011010010110011100100110010010000010011000101000010100010110000000110010010000110100100101011101001000110110100010110010110010001110000001111001101001110101000111000000001101111101011100101100001110101011110001001101100101011010010001000010101101001110000011100110011110100111001011111100010101110000101011010111000010010011100100001011110011001100100100011101101111100100101111110111101010011101010101001101001010101100100011010101111111111000011101110100110010111000000001000001110001001001010110000001010010000000111010111000010100101010101000010001010111000000101110111101100101000001000001000111111011011000011110010110111000111000000001111111011000000101111101011010111110111011111001110111100001011111111000000111111001101010101000000000001001000001100111010010011001000100010011011011111011100001111010001110010110111110101010101011100110000100001100111011000110100110110100100100011000011001100100111000010000100001000010101100001101011011100010111001010100100011100010111001000001010000101010111001111011110110001110101110000111101001010100010011010110100100101001000111001100010111101100101010110110110010100111111100110111000011110100011000101000110000001010111111011001011010111101000010100100010100110000001110010101010101010111001111010010111110001111010001101001010001011000101011100010001000001111010010101011100110100000010100001101110010100000010101001100010010011011110000000101001001011011100011000100101011110010101010101001010000001101011110011111011110110001011101001011011000100011001100110011111110111110010101011001100111111010010100011100011011010001010111110001111011001101010010001010101010010100001000110011100110000011111101000100110011011110110110011011001110110010010100110010100010110011011010100100000100010100100001000000011000111011011011100000100100110011010111010110001001111001010011110100101101111011001100110111000110011101011101010111101010000101111110011010000001001100011110011111011100010100001001001001000001100011000000111001111000111101101110011101010001111010011000111110011111100110001001010000000101010010100011111011010000110111111100000000011101111110010101111001000111111010000101000001010101101010000101101111011100001111111001100111101100001001111011001001010011111000011100001000011100110000000000111101000010011000110111111101001011001010100001011010011011011001110100000001000111100100001100110100100001101100101000101110010100111110111111001100010111011111111000011101110011001000011010001111100011100000001111000111110000010011111111111100101110010000111011011000000101010001100110000111101100001111111011001000011100100110000000011000100011000001100101110101101110110110001010010100000110011110011000111111001001000110000010100010011100010000011000010001100101101000101001111110101011111111101000101101001111000111111110110111010100000101100100100001111011110011110101010101011011100110110001110111011000101011010110111000000000001010110110001110000101001100001011010111010001101011011000000010000010000110111101101100000001111010100101101011011011100001100101001111000000010010011010010000001000111010001001010110000101010010100110111010110001101110001011110110010000100101111110010110011011100001010000000101010000001010000100011111111000001000011111010000100001100011011001100100000001000100110011110100110111000010000101100101000011011101010011000101100011110011111111100011100110110100110011111001001110000100001111100101011110001011010000010101001111111010001100000111100110110010110110010011101001001011000100000011010111101000001011000011001010001001001000101100000011100110000100000110101010;
wire[23:0] cb2_crc = 24'b001010100010111010110100;
wire[6143:0] output_vector2 = {cb2_crc, cb2_data};

//Clock Generator
initial clk=1'b0;
always #5 clk=~clk;


//Continously Readout the output buffer
always@(posedge clk, reset) begin
	if(reset==1'b1) begin
		rreq_itl <= 1'b0;
		rreq_enc <= 1'b0;
	end
	else begin
		if(empty_itl==1'b0)
			rreq_itl <= 1'b1;
		else
			rreq_itl <= 1'b0;
		
		if(empty_enc==1'b0)
			rreq_enc <= 1'b1;
		else
			rreq_enc <= 1'b0;
	end
end 


//Power-on Reset
initial
begin
		reset = 1'b1;
#20 	reset = 1'b0;
end


initial
begin	
	wreq_size = 1'b0;
	wreq_tb = 1'b0;
	tb_size_in = 16'b0;
	tb_in = 8'b0;
end

initial
begin
#50	wreq_size = 1'b1;
		tb_size_in = length;
#15	wreq_size = 1'b0;
#25	wreq_tb = 1'b1;
#5
	i = 0;
	k = -1;
	while (i < iterations)
	begin
		//#10 
		
		if (i < length) 
			tb_in = input_vector[i*8 +: 8];
		else
			tb_in = 0;
		
		//if (record_start == 1'b1 & k < 1056 & switch == 1'b0)
		if (record_start == 1'b1 & k < 132 & switch == 1'b0)
			begin
				if(k>-1)
					check_out = output_vector1[k*8 +: 8];
				k = k + 1;
			end
		//else if (record_start == 1'b1 &  k < 6144 & switch == 1'b1)
		else if (record_start == 1'b1 &  k < 768 & switch == 1'b1)
			begin
				if(k>-1)
					check_out = output_vector2[k*8 +: 8];
				k = k + 1;			
			end		
		else
			check_out = 0;
		i = i + 1;
		#10;
	end

end

initial 
begin

repeat(length * 20) 
	begin
	#1
		if (start_itl == 1'b1)
			begin
				record_start = 1'b1;
			end
		
		//if (record_start == 1'b1 & k==1056 & switch == 1'b0)
		if (record_start == 1'b1 & k==132 & switch == 1'b0)
			begin
				record_start = 1'b0;
				switch = 1'b1;
				k = -1;
			end
	end
end

endmodule
