`timescale 1ns/1ps
module tb_cb_seg();
reg clk, reset, tb_in, wreq_tb, wreq_size;

reg[15:0] tb_size_in;

wire empty_itl,empty_enc;
reg  rreq_itl, rreq_enc;

wire[2:0] q_enc;
wire data_enc, size_enc, start_enc;

wire[4:0] q_itl;
wire data_itl, size_itl, start_itl, crc_itl, filling_itl;


cb_seg test_obj(
    .clk(clk),
    .reset(reset),
    .tb_in(tb_in),
    .wreq_data(wreq_tb),
    .tb_size_in(tb_size_in),  
    .wreq_size(wreq_size),
	 
	 .rreq_itl_fifo(rreq_itl),
	 .q_itl_fifo(q_itl), //{data, size, start}
	 .empty_itl_fifo(empty_itl),
	 
	 //Encoder FIFO Ports
	 .rreq_enc_fifo(rreq_enc),
	 .q_enc_fifo(q_enc),  //{data, size, start, crc, filling}
	 .empty_enc_fifo(empty_enc)
	 
//
//    .filling(filling),
//    .crc(crc),
//    .start(start),
//    //.stop(stop),
//    .cb_size(cb_size),
//    .cb_data(cb_data) 
);

assign data_enc = q_enc[2];
assign size_enc = q_enc[1];
assign start_enc = q_enc[0];

assign data_itl = q_itl[4];
assign size_itl = q_itl[3];
assign start_itl = q_itl[2];
assign crc_itl = q_itl[1];
assign filling_itl = q_itl[0];

integer length = 7010;
integer iterations = 7250, i, k;
integer record_start= 0;
reg check_out, switch = 1'b0;

wire[7009:0] input_vector = 7010'b01010111010000111110001010010101011011111101101010101110000010110010001010010000111111001100011100010000100001101111000100101011010111100000011001011101100101101111101010011010111110011011000111011110010111000101101111001000111101001001101100111001000001111101001000000001000101001101101001001100000100111010000101110001100011011000111100010101101111111110110011100010111000101110001001110010101111010110100011000101010011011000001010011011001111110110011101100000111000111011111110100000011000100001001001001111011000010000101101010000010001110100011000111001100100001011000101010101000010101001101001001101011000010111010010011110010000010110010100010001111011000001010100100110100000100110011011011000111100111110000000000000110011001101001010101001001000100000101011110100100101111110100110001101000011011011000001001011100100101100001001101001101111100000010010111000010100000101010100011100111111101011111001011111110101110010110010101011010001110000001011111110100111011101011100000000011000111101010110111110000110010010001111000111110100010110010101111000000001000010001111101101010010011001100011000110111111111100110001011101100101101011111101001010110001101000101111110110011001000010000011011101101101100010111001101011100110010100001010111000000110011011110000100100100100011111011011100111000000011100000101010001000000001011001000000110111111001110011010000000101111011111010000010101110011111010101010110000110010101100000110101000100010110001110001110010001100011100011101100101100111001001110011001110000100011001001001010101110011101100000101000000100000100100111010010001110010011110000000101101100001010000011011001111010111001010001110111101000110101000011100000011111111010111010001111100001101101100101100101100010100011110101110010111000100100100100100111100001101011000100011011010001100010101101011000001111100010000000100100011011001101101111010111111110010000010111101001111001111101101111101001010011110001110110010110000011111110011100101111101111101101011011100000101100100101100011100011100101100101011110011001111001011000011011110100101110011010100111101111100000111111100101101101000101001111100101001000011010111011101010010011100001101110101111101111110001111000110000000110011001001110000011100010000110000111110110001010101001110111111000101111111110001010101001010101111011101011110011110101101000100000111011001011010010111111001100100101000001000011111111110110111000110000101110111010101100101001011001110001001011010001000111100101101101000111001001111111100011000010000111001010100110011000101010001011110110101101001011001110010011001001000001001100010100001010001011000000011001001000011010010010101110100100011011010001011001011001000111000000111100110100111010100011100000000110111110101110010110000111010101111000100110110010101101001000100001010110100111000001110011001111010011100101111110001010111000010101101011100001001001110010000101111001100110010010001110110111110010010111111011110101001110101010100110100101010110010001101010111111111100001110111010011001011100000000100000111000100100101011000000101001000000011101011100001010010101010100001000101011100000010111011110110010100000100000100011111101101100001111001011011100011100000000111111101100000010111110101101011111011101111100111011110000101111111100000011111100110101010100000000000100100000110011101001001100100010001001101101111101110000111101000111001011011111010101010101110011000010000110011101100011010011011010010010001100001100110010011100001000010000100001010110000110101101110001011100101010010001110001011100100000101000010101011100111101111011000111010111000011110100101010001001101011010010010100100011100110001011110110010101011011011001010011111110011011100001111010001100010100011000000101011111101100101101011110100001010010001010011000000111001010101010101011100111101001011111000111101000110100101000101100010101110001000100000111101001010101110011010000001010000110111001010000001010100110001001001101111000000010100100101101110001100010010101111001010101010100101000000110101111001111101111011000101110100101101100010001100110011001111111011111001010101100110011111101001010001110001101101000101011111000111101100110101001000101010101001010000100011001110011000001111110100010011001101111011011001101100111011001001010011001010001011001101101010010000010001010010000100000001100011101101101110000010010011001101011101011000100111100101001111010010110111101100110011011100011001110101110101011110101000010111111001101000000100110001111001111101110001010000100100100100000110001100000011100111100011110110111001110101000111101001100011111001111110011000100101000000010101001010001111101101000011011111110000000001110111111001010111100100011111101000010100000101010110101000010110111101110000111111100110011110110000100111101100100101001111100001110000100001110011000000000011110100001001100011011111110100101100101010000101101001101101100111010000000100011110010000110011010010000110110010100010111001010011111011111100110001011101111111100001110111001100100001101000111110001110000000111100011111000001001111111111110010111001000011101101100000010101000110011000011110110000111111101100100001110010011000000001100010001100000110010111010110111011011000101001010000011001111001100011111100100100011000001010001001110001000001100001000110010110100010100111111010101111111110100010110100111100011111111011011101010000010110010010000111101111001111010101010101101110011011000111011101100010101101011011100000000000101011011000111000010100110000101101011101000110101101100000001000001000011011110110110000000111101010010110101101101110000110010100111100000001001001101001000000100011101000100101011000010101001010011011101011000110111000101111011001000010010111111001011001101110000101000000010101000000101000010001111111100000100001111101000010000110001101100110010000000100010011001111010011011100001000010110010100001101110101001100010110001111001111111110001110011011010011001111100100111000010000111110010101111000101101000001010100111111101000110000011110011011001011011001001110100100101100010000001101011110100000101100001100101000100100100010110000001110011000010000011010101011110110100010101111001110110111101101111100000100010001111111110000000100011000011110101111111000011000111101110100111000011000110101001100110011110001001010001110000111001100101010110000110110000000000000101001001000111111111100010000101111000001110001000100101101000001011100110101101001010110110001111110001110110110000100011010100010100100010111111110011000010000100011100011111101011110110111011011101011110000101011001111111110010001000101000000100000100001000010111100100101001110110110100111000111001000000110110100010010110010011110101110001111000010000101100101011011100011100010011001101111100011100111001001111001100000011001001100100101011100000000110100011001001010111101010101111001111011011111001001110001001011111100010000010111010001010010011001011011010101001001001001000000010010101110110011010101111000100100100000000100000111010100101011010111100010010111001111101110;

wire[1031:0] cb1_data = 1032'b111101101000101011110011101101111011011111000001000100011111111100000001000110000111101011111110000110001111011101001110000110001101010011001100111100010010100011100001110011001010101100001101100000000000001010010010001111111111000100001011110000011100010001001011010000010111001101011010010101101100011111100011101101100001000110101000101001000101111111100110000100001000111000111111010111101101110110111010111100001010110011111111100100010001010000001000001000010000101111001001010011101101101001110001110010000001101101000100101100100111101011100011110000100001011001010110111000111000100110011011111000111001110010011110011000000110010011001001010111000000001101000110010010101111010101011110011110110111110010011100010010111111000100000101110100010100100110010110110101010010010010010000000100101011101100110101011110001001001000000001000001110101001010110101111000100101110011111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire[23:0] cb1_crc = 24'b011110101001100101000010;
//From MSB to LSB
wire[1055:0] output_vector1 = {cb1_crc, cb1_data};


wire[6119:0] cb2_data = 6120'b010101110100001111100010100101010110111111011010101011100000101100100010100100001111110011000111000100001000011011110001001010110101111000000110010111011001011011111010100110101111100110110001110111100101110001011011110010001111010010011011001110010000011111010010000000010001010011011010010011000001001110100001011100011000110110001111000101011011111111101100111000101110001011100010011100101011110101101000110001010100110110000010100110110011111101100111011000001110001110111111101000000110001000010010010011110110000100001011010100000100011101000110001110011001000010110001010101010000101010011010010011010110000101110100100111100100000101100101000100011110110000010101001001101000001001100110110110001111001111100000000000001100110011010010101010010010001000001010111101001001011111101001100011010000110110110000010010111001001011000010011010011011111000000100101110000101000001010101000111001111111010111110010111111101011100101100101010110100011100000010111111101001110111010111000000000110001111010101101111100001100100100011110001111101000101100101011110000000010000100011111011010100100110011000110001101111111111001100010111011001011010111111010010101100011010001011111101100110010000100000110111011011011000101110011010111001100101000010101110000001100110111100001001001001000111110110111001110000000111000001010100010000000010110010000001101111110011100110100000001011110111110100000101011100111110101010101100001100101011000001101010001000101100011100011100100011000111000111011001011001110010011100110011100001000110010010010101011100111011000001010000001000001001001110100100011100100111100000001011011000010100000110110011110101110010100011101111010001101010000111000000111111110101110100011111000011011011001011001011000101000111101011100101110001001001001001001111000011010110001000110110100011000101011010110000011111000100000001001000110110011011011110101111111100100000101111010011110011111011011111010010100111100011101100101100000111111100111001011111011111011010110111000001011001001011000111000111001011001010111100110011110010110000110111101001011100110101001111011111000001111111001011011010001010011111001010010000110101110111010100100111000011011101011111011111100011110001100000001100110010011100000111000100001100001111101100010101010011101111110001011111111100010101010010101011110111010111100111101011010001000001110110010110100101111110011001001010000010000111111111101101110001100001011101110101011001010010110011100010010110100010001111001011011010001110010011111111000110000100001110010101001100110001010100010111101101011010010110011100100110010010000010011000101000010100010110000000110010010000110100100101011101001000110110100010110010110010001110000001111001101001110101000111000000001101111101011100101100001110101011110001001101100101011010010001000010101101001110000011100110011110100111001011111100010101110000101011010111000010010011100100001011110011001100100100011101101111100100101111110111101010011101010101001101001010101100100011010101111111111000011101110100110010111000000001000001110001001001010110000001010010000000111010111000010100101010101000010001010111000000101110111101100101000001000001000111111011011000011110010110111000111000000001111111011000000101111101011010111110111011111001110111100001011111111000000111111001101010101000000000001001000001100111010010011001000100010011011011111011100001111010001110010110111110101010101011100110000100001100111011000110100110110100100100011000011001100100111000010000100001000010101100001101011011100010111001010100100011100010111001000001010000101010111001111011110110001110101110000111101001010100010011010110100100101001000111001100010111101100101010110110110010100111111100110111000011110100011000101000110000001010111111011001011010111101000010100100010100110000001110010101010101010111001111010010111110001111010001101001010001011000101011100010001000001111010010101011100110100000010100001101110010100000010101001100010010011011110000000101001001011011100011000100101011110010101010101001010000001101011110011111011110110001011101001011011000100011001100110011111110111110010101011001100111111010010100011100011011010001010111110001111011001101010010001010101010010100001000110011100110000011111101000100110011011110110110011011001110110010010100110010100010110011011010100100000100010100100001000000011000111011011011100000100100110011010111010110001001111001010011110100101101111011001100110111000110011101011101010111101010000101111110011010000001001100011110011111011100010100001001001001000001100011000000111001111000111101101110011101010001111010011000111110011111100110001001010000000101010010100011111011010000110111111100000000011101111110010101111001000111111010000101000001010101101010000101101111011100001111111001100111101100001001111011001001010011111000011100001000011100110000000000111101000010011000110111111101001011001010100001011010011011011001110100000001000111100100001100110100100001101100101000101110010100111110111111001100010111011111111000011101110011001000011010001111100011100000001111000111110000010011111111111100101110010000111011011000000101010001100110000111101100001111111011001000011100100110000000011000100011000001100101110101101110110110001010010100000110011110011000111111001001000110000010100010011100010000011000010001100101101000101001111110101011111111101000101101001111000111111110110111010100000101100100100001111011110011110101010101011011100110110001110111011000101011010110111000000000001010110110001110000101001100001011010111010001101011011000000010000010000110111101101100000001111010100101101011011011100001100101001111000000010010011010010000001000111010001001010110000101010010100110111010110001101110001011110110010000100101111110010110011011100001010000000101010000001010000100011111111000001000011111010000100001100011011001100100000001000100110011110100110111000010000101100101000011011101010011000101100011110011111111100011100110110100110011111001001110000100001111100101011110001011010000010101001111111010001100000111100110110010110110010011101001001011000100000011010111101000001011000011001010001001001000101100000011100110000100000110101010;
wire[23:0] cb2_crc = 24'b001010100010111010110100;
wire[6143:0] output_vector2 = {cb2_crc, cb2_data};

//Clock Generator
initial clk=1'b0;
always #5 clk=~clk;


//Continously Readout the output buffer
always@(posedge clk, reset) begin
	if(reset==1'b1) begin
		rreq_itl <= 1'b0;
		rreq_enc <= 1'b0;
	end
	else begin
		if(empty_itl==1'b0)
			rreq_itl <= 1'b1;
		else
			rreq_itl <= 1'b0;
		
		if(empty_enc==1'b0)
			rreq_enc <= 1'b1;
		else
			rreq_enc <= 1'b0;
	end
end 


//Power-on Reset
initial
begin
		reset = 1'b1;
#20 	reset = 1'b0;
end


initial
begin	
	wreq_size = 1'b0;
	wreq_tb = 1'b0;
	tb_size_in = 16'h0;
	tb_in = 1'b0;
end

initial
begin
#50	wreq_size = 1'b1;
		tb_size_in = length;
#15	wreq_size = 1'b0;
#25	wreq_tb = 1'b1;
#5
	i = 0;
	k = -1;
	while (i < iterations)
	begin
		//#10 
		
		if (i < 7010) 
			tb_in = input_vector[i];
		else
			tb_in = 0;
		
		if (record_start == 1'b1 & k < 1056 & switch == 1'b0)
			begin
				if(k>-1)
					check_out = output_vector1[k];
				k = k + 1;
			end
		else if (record_start == 1'b1 &  k < 6144 & switch == 1'b1)
			begin
				if(k>-1)
					check_out = output_vector2[k];
				k = k + 1;			
			end		
		else
			check_out = 0;
		i = i + 1;
		#10;
	end

end

initial 
begin

repeat(length * 20) 
	begin
	#1
		if (start_itl == 1'b1)
			begin
				record_start = 1'b1;
			end
		
		if (record_start == 1'b1 & k==1056 & switch == 1'b0)
			begin
				record_start = 1'b0;
				switch = 1'b1;
				k = -1;
			end
	end
end

endmodule
