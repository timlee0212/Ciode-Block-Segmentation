//`timescale 1ns/1ps
//module tb_control_path();
//
//reg clk, reset;
//
//always #5 clk = ~clk;  //100MHz
//
//initial
//begin
//	reset = 1'b1;
//	#20
//	
//end
//
//endmodule